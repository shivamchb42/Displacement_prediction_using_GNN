b0VIM 8.2      YH c�
 G1  piyush                                  piyush-Latitude-3460                    ~piyush/Documents/piyushFEM/femcode2 (4) _fgm/cont_ver2/shape                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      3210    #"! U                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 tp           g                                   h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      ad     �     g       �  �  �  �  �  �  7      �  �  �  �    |  G      �  �  �  �  |  V  0  
  �  �  �  �  [  /    �  �    S  '  �
  �
  �
  �
  �
  �
  m
  I
  %
  
  �	  �	  �	  q	  [	  >	  	  �  �  �  |  P  $  �  �  �  t  H    �  �  �  �  x  g  C    �  �  �  �  k  G  #    �  �  �  �  �  I  F  4  (  &    �  �  M    �  �  M    �  �                        displacement 9  2.105044978349781E-010 -7.464602743625567E-012  displacement 8  2.284915845212138E-010  7.492285333427082E-026  displacement 7  2.105044978349781E-010  7.464602743625693E-012  displacement 6  1.447925255924183E-010 -3.245823406756952E-011  displacement 5  1.478367889782390E-010  3.231174267785264E-026  displacement 4  1.447925255924185E-010  3.245823406756959E-011  displacement 3  0.000000000000000E+000  0.000000000000000E+000  displacement 2  0.000000000000000E+000  0.000000000000000E+000  displacement 1  0.000000000000000E+000  0.000000000000000E+000   0.000000000000000E+000    hybpr ends  cint           2     ratnorm = |{unbal}|/|{f_incr}| =  0.1732E-09 < equitol    sqn_unbal,sqn_ldtdt   0.5398E-16  0.1800E+04   1.000000000000000E-008  sum glbld -    60.0000000000000       time in elem  1.9999999E-04   Subroutine stiffp99  x0 in celt   1.00000000000000       x0 in celt  0.225403330758517       x0 in celt   1.00000000000000       x0 in celt   1.77459666924148       x0 in celt   1.00000000000000       x0 in celt  0.225403330758517       x0 in celt   1.77459666924148       x0 in celt   1.77459666924148       x0 in celt  0.225403330758517      .. Iteration   2 .. Factor   0.1000000E+01    1      1.00000000000000                1  3.3820000E-02  0.1361710      up9  3.3299625E-04  x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds  0.225403330758517       x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds  0.225403330758517       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds  0.225403330758517       berr  5.329070518200751E-016  ratnorm = |{unbal}|/|{f_incr}| =  0.1000E+01 > equitol sqn_unbal,sqn_ldtdt   0.1800E+04  0.1800E+04   1.000000000000000E-008  sum glbld -    60.0000000000000       time in elem  3.0000001E-04   Subroutine stiffp99  x0 in celt   1.00000000000000       x0 in celt  0.225403330758517       x0 in celt   1.00000000000000       x0 in celt   1.77459666924148       x0 in celt   1.00000000000000       x0 in celt  0.225403330758517       x0 in celt   1.77459666924148       x0 in celt   1.77459666924148       x0 in celt  0.225403330758517      .. Iteration   1 .. Factor   0.1000000E+01    1    up9  3.5000220E-04  x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds  0.225403330758517       x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds   1.00000000000000       x0 in upaspeloi2ds  0.225403330758517       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds   1.77459666924148       x0 in upaspeloi2ds  0.225403330758517       iarc, ichord            0           1  nmvalues          144   Number of equations =           12   > ... Input data is complete.   >> ... User-typed input is complete   >> ... User-typed input is complete   >> ... User-typed input is complete   >> ... User-typed input is complete  contfc2 -   contfc1 -   end of contread   0.000000000000000E+000  0.000000000000000E+000  0.000000000000000E+000      0 0.100E+01 0.100E+01     0     0     0     1  mflg2,maxtime,deltat , ipress,igrav,icont,loadsteps     in contread  You can modify the parameter mx_incdim to            9  cl -            1 ,clsspt -           1  in eledefi  p9_3                  0           0            1           9  Analysis for,q4 combined geometry  9  nodes   1    elements                       >>> Subroutine ctrldata  plane stress   Restart program using a data file ?        Subroutine intarray   Program main ad  �  �            �  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                ********************************* 